library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;
  use IEEE.std_logic_unsigned.all;

entity NOMBRE is
  port (entrada1 : in  std_logic;
        entrada2 : in  std_logic_vector(4 downto 0);
        salida1  : out std_logic;
        salida2  : out std_logic_vector(5 downto 0)
       );
end entity;

architecture Behavioral of NOMBRE is
  -- COMPONENTS SIGNALS
begin
  --DISENO
end architecture;

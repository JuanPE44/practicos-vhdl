library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;
  use IEEE.std_logic_unsigned.all;

entity NOMBRE is
  port (entrada1 : in  STD_LOGIC;
        entrada2 : in  STD_LOGIC_VECTOR(4 downto 0);
        salida1  : out STD_LOGIC;
        salida2  : out STD_LOGIC_VECTOR(5 downto 0)
       );
end entity;

architecture Behavioral of NOMBRE is
  -- COMPONENTS SIGNALS
begin
  --DISENO
end architecture;
